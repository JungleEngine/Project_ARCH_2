LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DECODER IS
	Port ( 
		X : IN STD_LOGIC_VECTOR (2 downto 0);
	  EN : IN std_logic;
		Y : OUT STD_LOGIC_VECTOR (5 downto 0)
		);
END DECODER;

ARCHITECTURE BEHAVIORAL OF DECODER IS
BEGIN
	     Y <= "000001" WHEN (X = "000" AND EN = '1')
	     ELSE "000010" WHEN (X = "001" AND EN = '1')
	     ELSE "000100" WHEN (X = "010" AND EN = '1')
	     ELSE "001000" WHEN (X = "011" AND EN = '1')
	     ELSE "010000" WHEN (X = "100" AND EN = '1')
	     ELSE "100000" WHEN (X = "101" AND EN = '1')
	     ELSE "000000";
END BEHAVIORAL;