LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;
USE IEEE.STD_LOGIC_SIGNED.all;

ENTITY REG_FILE IS
	GENERIC(N : integer := 16);
		PORT(
			CLK: IN std_logic;
			RST: IN std_logic;

			SP_INC: IN std_logic;
			SP_DEC: IN std_logic;
			PC_ENABLE: IN std_logic;
			WB_FR_ENABLE: IN std_logic;
			ALU_FR_ENABLE: IN std_logic;
			DECODE_FR_ENABLE: IN std_logic;

			WB_Rdst_INDEX: IN std_logic_vector(2 downto 0);
			WB_Rsrc_INDEX: IN std_logic_vector(2 downto 0);
			ALU_Rdst_INDEX: IN std_logic_vector(2 downto 0);
			ALU_Rsrc_INDEX: IN std_logic_vector(2 downto 0);
			DECODE_Rdst_INDEX: IN std_logic_vector(2 downto 0);

			PC_IN_DATA: IN std_logic_vector(8 DOWNTO 0);
			WB_FR_DATA: IN std_logic_vector(3 DOWNTO 0);
			ALU_FR_DATA: IN std_logic_vector(3 DOWNTO 0);
			DECODE_FR_DATA: IN std_logic_vector(3 DOWNTO 0);
			IN_BUS: IN std_logic_vector(31 DOWNTO 0);

			ALU_OUT_BUS: OUT std_logic_vector(31 DOWNTO 0);
			DECODE_OUT_BUS: OUT std_logic_vector(15 DOWNTO 0);

			PC_OUT_DATA: OUT std_logic_vector(8 DOWNTO 0);
			SP_OUT_DATA: OUT std_logic_vector(8 DOWNTO 0);
			FR_OUT_DATA: OUT std_logic_vector(3 DOWNTO 0)
		);
END REG_FILE;

ARCHITECTURE REG_FILE_ARCH OF REG_FILE IS

SIGNAL SP_VALUE: std_logic_vector(8 DOWNTO 0);
SIGNAL R0_IN_DATA: std_logic_vector(15 DOWNTO 0);
SIGNAL R1_IN_DATA: std_logic_vector(15 DOWNTO 0);
SIGNAL R2_IN_DATA: std_logic_vector(15 DOWNTO 0);
SIGNAL R3_IN_DATA: std_logic_vector(15 DOWNTO 0);
SIGNAL R4_IN_DATA: std_logic_vector(15 DOWNTO 0);
SIGNAL R5_IN_DATA: std_logic_vector(15 DOWNTO 0);
SIGNAL FR_IN_DATA: std_logic_vector(3 DOWNTO 0);
SIGNAL SP_IN_DATA: std_logic_vector(8 DOWNTO 0);

SIGNAL R0_OUT_DATA: std_logic_vector(15 DOWNTO 0);
SIGNAL R1_OUT_DATA: std_logic_vector(15 DOWNTO 0);
SIGNAL R2_OUT_DATA: std_logic_vector(15 DOWNTO 0);
SIGNAL R3_OUT_DATA: std_logic_vector(15 DOWNTO 0);
SIGNAL R4_OUT_DATA: std_logic_vector(15 DOWNTO 0);
SIGNAL R5_OUT_DATA: std_logic_vector(15 DOWNTO 0);

SIGNAL FR_ENABLE: std_logic;
SIGNAL SP_ENABLE: std_logic;
SIGNAL R0_ENABLE: std_logic;
SIGNAL R1_ENABLE: std_logic;
SIGNAL R2_ENABLE: std_logic;
SIGNAL R3_ENABLE: std_logic;
SIGNAL R4_ENABLE: std_logic;
SIGNAL R5_ENABLE: std_logic;
SIGNAL WB_REGISTERS_WRITE_ENABLES_LSB: std_logic_vector(5 DOWNTO 0);
SIGNAL WB_REGISTERS_WRITE_ENABLES_MSB: std_logic_vector(5 DOWNTO 0);
SIGNAL ALU_REGISTERS_WRITE_ENABLES_LSB: std_logic_vector(5 DOWNTO 0);
SIGNAL ALU_REGISTERS_WRITE_ENABLES_MSB: std_logic_vector(5 DOWNTO 0);
SIGNAL DECODE_REGISTERS_WRITE_ENABLES: std_logic_vector(5 DOWNTO 0);
SIGNAL NOT_CLK: std_logic;

BEGIN
	
	NOT_CLK<= not CLK;
	
	SP_ENABLE <= '1' WHEN (SP_DEC = '1' AND SP_INC = '0') OR (SP_INC = '1' AND SP_DEC = '0')
	ELSE '0';

	FR_ENABLE <= '1'  WHEN (WB_FR_ENABLE = '1' OR DECODE_FR_ENABLE = '1' OR ALU_FR_ENABLE = '1')
	ELSE '0';

	R0_ENABLE <= '1' WHEN WB_REGISTERS_WRITE_ENABLES_LSB(0) = '1' or WB_REGISTERS_WRITE_ENABLES_MSB(0) = '1'
	ELSE '0';

	R1_ENABLE <= '1' WHEN WB_REGISTERS_WRITE_ENABLES_LSB(1) = '1' or WB_REGISTERS_WRITE_ENABLES_MSB(1) = '1'
	ELSE '0';

	R2_ENABLE <= '1' WHEN WB_REGISTERS_WRITE_ENABLES_LSB(2) = '1' or WB_REGISTERS_WRITE_ENABLES_MSB(2) = '1'
	ELSE '0';

	R3_ENABLE <= '1' WHEN WB_REGISTERS_WRITE_ENABLES_LSB(3) = '1' or WB_REGISTERS_WRITE_ENABLES_MSB(3) = '1'
	ELSE '0';

	R4_ENABLE <= '1' WHEN WB_REGISTERS_WRITE_ENABLES_LSB(4) = '1' or WB_REGISTERS_WRITE_ENABLES_MSB(4) = '1'
	ELSE '0';

	R5_ENABLE <= '1' WHEN WB_REGISTERS_WRITE_ENABLES_LSB(5) = '1' or WB_REGISTERS_WRITE_ENABLES_MSB(5) = '1'
	ELSE '0';


  SP_OUT_DATA <= SP_VALUE;
  
	SP_IN_DATA <= (SP_VALUE + 1) WHEN (SP_INC = '1')
	ELSE (SP_VALUE - 1) WHEN (SP_DEC = '1')
	ELSE SP_VALUE;

	FR_IN_DATA <= WB_FR_DATA WHEN (WB_FR_ENABLE = '1')
	ELSE DECODE_FR_DATA WHEN (DECODE_FR_ENABLE = '1')
	ELSE ALU_FR_DATA;
	  
	R0_IN_DATA <= IN_BUS(15 DOWNTO 0) WHEN WB_REGISTERS_WRITE_ENABLES_LSB(0) = '1'
	ELSE IN_BUS(31 DOWNTO 16);

	R1_IN_DATA <= IN_BUS(15 DOWNTO 0) WHEN WB_REGISTERS_WRITE_ENABLES_LSB(1) = '1'
	ELSE IN_BUS(31 DOWNTO 16);

	R2_IN_DATA <= IN_BUS(15 DOWNTO 0) WHEN WB_REGISTERS_WRITE_ENABLES_LSB(2) = '1'
	ELSE IN_BUS(31 DOWNTO 16);

	R3_IN_DATA <= IN_BUS(15 DOWNTO 0) WHEN WB_REGISTERS_WRITE_ENABLES_LSB(3) = '1'
	ELSE IN_BUS(31 DOWNTO 16);

	R4_IN_DATA <= IN_BUS(15 DOWNTO 0) WHEN WB_REGISTERS_WRITE_ENABLES_LSB(4) = '1'
	ELSE IN_BUS(31 DOWNTO 16);

	R5_IN_DATA <= IN_BUS(15 DOWNTO 0) WHEN WB_REGISTERS_WRITE_ENABLES_LSB(5) = '1'
	ELSE IN_BUS(31 DOWNTO 16);


	ALU_OUT_BUS(15 DOWNTO 0) <= R0_OUT_DATA WHEN ALU_REGISTERS_WRITE_ENABLES_LSB(0) = '1'
	ELSE R1_OUT_DATA WHEN ALU_REGISTERS_WRITE_ENABLES_LSB(1) = '1'
	ELSE R2_OUT_DATA WHEN ALU_REGISTERS_WRITE_ENABLES_LSB(2) = '1'
	ELSE R3_OUT_DATA WHEN ALU_REGISTERS_WRITE_ENABLES_LSB(3) = '1'
	ELSE R4_OUT_DATA WHEN ALU_REGISTERS_WRITE_ENABLES_LSB(4) = '1'
	ELSE R5_OUT_DATA WHEN ALU_REGISTERS_WRITE_ENABLES_LSB(5) = '1';


	ALU_OUT_BUS(31 DOWNTO 16) <= R0_OUT_DATA WHEN ALU_REGISTERS_WRITE_ENABLES_MSB(0) = '1'
	ELSE R1_OUT_DATA WHEN ALU_REGISTERS_WRITE_ENABLES_MSB(1) = '1'
	ELSE R2_OUT_DATA WHEN ALU_REGISTERS_WRITE_ENABLES_MSB(2) = '1'
	ELSE R3_OUT_DATA WHEN ALU_REGISTERS_WRITE_ENABLES_MSB(3) = '1'
	ELSE R4_OUT_DATA WHEN ALU_REGISTERS_WRITE_ENABLES_MSB(4) = '1'
	ELSE R5_OUT_DATA WHEN ALU_REGISTERS_WRITE_ENABLES_MSB(5) = '1';


	DECODE_OUT_BUS <= R0_OUT_DATA WHEN DECODE_REGISTERS_WRITE_ENABLES(0) = '1'
	ELSE R1_OUT_DATA WHEN DECODE_REGISTERS_WRITE_ENABLES(1) = '1'
	ELSE R2_OUT_DATA WHEN DECODE_REGISTERS_WRITE_ENABLES(2) = '1'
	ELSE R3_OUT_DATA WHEN DECODE_REGISTERS_WRITE_ENABLES(3) = '1'
	ELSE R4_OUT_DATA WHEN DECODE_REGISTERS_WRITE_ENABLES(4) = '1'
	ELSE R5_OUT_DATA WHEN DECODE_REGISTERS_WRITE_ENABLES(5) = '1';

	-- Decoder to generate register enable signals from Rsrc and Rdst indexes
	WB_REGISTERS_DECODER_LSB: ENTITY work.DECODER PORT MAP (WB_Rsrc_INDEX, WB_REGISTERS_WRITE_ENABLES_MSB);
	WB_REGISTERS_DECODER_MSB: ENTITY work.DECODER PORT MAP (WB_Rdst_INDEX, WB_REGISTERS_WRITE_ENABLES_LSB);
	ALU_REGISTERS_DECODER_LSB: ENTITY work.DECODER PORT MAP (ALU_Rsrc_INDEX, ALU_REGISTERS_WRITE_ENABLES_LSB);
	ALU_REGISTERS_DECODER_MSB: ENTITY work.DECODER PORT MAP (ALU_Rdst_INDEX, ALU_REGISTERS_WRITE_ENABLES_MSB);
	DECODE_REGISTERS_DECODER_MSB: ENTITY work.DECODER PORT MAP (DECODE_Rdst_INDEX, DECODE_REGISTERS_WRITE_ENABLES);


	R0: ENTITY work.REG GENERIC MAP(n => 16) PORT MAP (R0_IN_DATA, R0_ENABLE,NOT_CLK, RST, R0_OUT_DATA);
	R1: ENTITY work.REG GENERIC MAP(n => 16) PORT MAP (R1_IN_DATA, R1_ENABLE, NOT_CLK, RST, R1_OUT_DATA);
	R2: ENTITY work.REG GENERIC MAP(n => 16) PORT MAP (R2_IN_DATA, R2_ENABLE, NOT_CLK, RST, R2_OUT_DATA);
	R3: ENTITY work.REG GENERIC MAP(n => 16) PORT MAP (R3_IN_DATA, R3_ENABLE, NOT_CLK, RST, R3_OUT_DATA);
	R4: ENTITY work.REG GENERIC MAP(n => 16) PORT MAP (R4_IN_DATA, R4_ENABLE, NOT_CLK, RST, R4_OUT_DATA);
	R5: ENTITY work.REG GENERIC MAP(n => 16) PORT MAP (R5_IN_DATA, R5_ENABLE, NOT_CLK, RST, R5_OUT_DATA);
	
	PC: ENTITY work.REG GENERIC MAP(n => 9) PORT MAP (PC_IN_DATA, PC_ENABLE, CLK, RST, PC_OUT_DATA);
	SP: ENTITY work.REG GENERIC MAP(n => 9) PORT MAP (SP_IN_DATA, SP_ENABLE, CLK, RST, SP_VALUE);
	FR: ENTITY work.REG GENERIC MAP(n => 4) PORT MAP (FR_IN_DATA, FR_ENABLE, CLK, RST, FR_OUT_DATA);


END REG_FILE_ARCH;